//!topmodule mkSimpleTest
module mkSimpleTest(Empty);
    
endmodule
