interface SecondModule;
endinterface

module mkSecondModule(SecondModule);
    method Bool isSecondModuleHookedUp;
        return True;
    endmethod
endmodule
