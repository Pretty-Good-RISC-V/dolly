//!topmodule mkSimpleTest
import Simple::*;

module mkSimpleTest(Empty);
    Simple simple <- mkSimple;
endmodule
