//!submodule embedded_module
