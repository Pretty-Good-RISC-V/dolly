//!submodule another_module
//!submodule second_module
